------------------------------------------------------------------------------------------------------------------------------------------
-- Project: Defender (DSD Final Project Fall 2021)
-- Author: Blake Martin & Nathan Gardner
-- Date: 11/30/21
------------------------------------------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package graphicsPackage is

	type point_2D is
	record
		x : integer;
		y : integer;
	end record;

	--CONSTANTS:
	constant mapEdgeLeft : integer := 0; -- leftmost pixel
	constant mapEdgeRight: integer := 640;
	constant mapEdgeTop :  integer := 30;
	constant mapEdgeBottom:integer := 460;
	constant COLS : integer := 640; --m
	constant ROWS : integer := 480;

    constant init_shipVel : integer := 0;
	constant shipsInitialx : integer := 150;
	constant shipsInitialy : integer := 240;

	--Ship geometry:
	constant shipHeightConst : integer := 25;
	constant shipWidthConst  : integer := 25;

    --Laser Geometry:
	constant laserWidth : integer := 10;
	constant laserHeight : integer := 2;

	-- enemy geometry
	constant smallHeight : integer := 15;
	constant smallWidth : integer  := 15;
	constant smallPoints : integer := 20;

	constant medHeight : integer := 25;
	constant medWidth : integer  := 25;
	constant medPoints : integer := 15;

	constant bigHeight : integer := 30;
	constant bigWidth : integer :=  30;
	constant bigPoints : integer := 10;
    --Enemey initial positions:
	constant smallStartX : integer := 645;
	constant smallStartY : integer := 100;
	constant medstartx   : integer := 645;
	constant medStartY   : integer := 350;
	constant bigStartX   : integer := 645;
	constant bigStartY   : integer := 300;

	constant objectWidth	 : integer := 25;
	constant objectHeight   : integer := 25;
	constant objPosX     : integer := 645;
	constant objPosy1     : integer := 212;
	constant objPosy2     : integer := 100;
	constant objPosy3     : integer := 420;
	constant objPosy4     : integer := 300;
	constant objPosy5     : integer := 150;
	constant objVeloX 	 : integer := -3;
	constant objVeloY    : integer := 0;
	--------------------------------------------------------------------------------------

	------ terrain --------------------added by Nathan-------------

	type terrain_type is array (1 to 10000) of integer;
		constant terrain_rom_const : terrain_type :=
		(
			1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,22,22,22,21,20,23,24,25,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,44,43,42,41,40,39,38,37,36,35,34,33,32,32,32,32,32,31,31,31,30,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0,1,2,3,4,5,6,7,8,9,10
		);
	type terrain_data is
		record
			pixelOn : boolean;
			rgb : std_logic_vector(11 downto 0);
		end record;
	constant init_terrain : terrain_data := (pixelOn => false, rgb => "011000110011");


	-----------------------------------------------------------------

--------------------- EXPLOSIONS ROMS -------------------------------------------------------------------------------------------------

	constant init_explosion_pos : point_2D := (x => 0, y => 0);

	type type_explosion is
	record
		position : point_2D;
		size : integer;
		pixelOn : boolean;
		rgb : std_logic_vector(11 downto 0);
		explosionHold : boolean;
	end record;
	constant init_explosion : type_explosion := (init_explosion_pos, 0, false, "111111111111", false);--- ****** ---

	type small_exp_rom_type is array (0 to 14) of std_logic_vector(0 to 14);
	constant small_exp_rom_const : small_exp_rom_type :=
	(
		"000000000000000",
		"000000100000000",
		"000000100010000",
		"000110111110000",
		"001011111111110",
		"111110000111110",
		"001100000001111",
		"111000000001111",
		"011100000001100",
		"011111000011111",
		"011011101111100",
		"000011111011000",
		"000010101000000",
		"000000001000000",
		"000000000000000"
	);

	type medium_exp_rom_type is array (0 to 24) of std_logic_vector(0 to 24);
	constant medium_exp_rom_const : medium_exp_rom_type :=
	(
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000100000000000000",
		"0000000000110000010000000",
		"0000110000110000110000000",
		"0000011000110110110000000",
		"0000001110101111100000110",
		"0000001111101010100111000",
		"1100111100100000111110000",
		"0111111110000000001101100",
		"0001100000000000001111000",
		"0000110000000000000111111",
		"0111100000000000000111100",
		"1111111000000000000110000",
		"0000110000000000000011000",
		"0011111010000000001111110",
		"0000111110000010011100011",
		"0001100010100011101111000",
		"0010000111111010111000000",
		"0000000110011110001100000",
		"0000000110010110000010000",
		"0000000100000110000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000"
	);


	type large_exp_rom_type is array (0 to 29) of std_logic_vector(0 to 29);
	constant large_exp_rom_const : large_exp_rom_type :=
	(
		"000000000000000000000000000000",
		"000000000000000000000000000000",
		"000000000000010000000000000000",
		"000000000000010000000100000000",
		"000000000000110000001100000000",
		"000001100000111010001100000000",
		"000000110000111010011000000000",
		"000000011100101111101000000110",
		"000000011110100111011000111100",
		"000011001001100000011111110000",
		"111101111100000000011001100000",
		"001111110100000000000011111100",
		"000111000000000000000111110000",
		"000001110000000000000001111111",
		"000111100000000000000000011111",
		"111100000000000000000011110000",
		"111111110000000000000001100000",
		"000001100000000000000000011000",
		"000111110010000000000011111110",
		"000000111110000001001111000111",
		"000011100110100001100111100000",
		"001110000101111101011010010000",
		"000000000101011111001110000000",
		"000000000110011110000011000000",
		"000000001100010010000001100000",
		"000000001000010010000000000000",
		"000000001000000010000000000000",
		"000000000000000000000000000000",
		"000000000000000000000000000000",
		"000000000000000000000000000000"
	);

-----------------------------------------------------------------------------

----------------------- MUSICAL NOTES FOR COUNTER ---------------------------

constant Asharp4 : std_logic_vector(23 downto 0) := "000000001000110010100010";
constant Dsharp4 : std_logic_vector(23 downto 0) := "000000001101001010111001";
constant Fsharp4 : std_logic_vector(23 downto 0) := "000000001011000100011111";


-----------------------------------------------------------------------------


	--NATHAN SCOREDBOARD / ROM UPDATES
	-- Variables related to the ROM for the ship ------------
	type rom_type is array (0 to 24) of std_logic_vector(0 to 24);
	constant ship_rom_const : rom_type :=
	(
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000011110000000000000000",
		"0000111110000000000000000",
		"0001111111000000000000000",
		"0001111111100000000000000",
		"0001111111111111111110000",
		"0001111111111111111111100",
		"0001111111111111111111110",
		"0000001111111000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000"
	);

	--- ship left and right boundry
	signal ship_x_l , ship_x_r : integer;
	--- ship top and bottom boundry
	signal ship_y_t , ship_y_b : integer;

	signal sq_ship_on : std_logic;

	signal ship_rom_addr , ship_rom_col : integer;
	signal ship_rom_data: std_logic_vector (0 to 24);
	signal ship_rom_bit : std_logic ;


------ Character set ROM --------------------------------------
-----------------------------------------------------------------

------ Variables related to the scoreboard ----------------------


	type scoreboard_data is
	record
		pixelOn : boolean;
		rgb : std_logic_vector(11 downto 0);
	end record;
	constant init_scoreboard : scoreboard_data := (pixelOn => false, rgb => "111001000011");

	type score_char is--- ****** ---
	record
		score_rom_opcode : std_logic_vector(6 downto 0);
		score_top : integer;
		score_bottom : integer;
		score_left : integer;
		score_right : integer;
		fontBitEn : std_logic;
		inScoreboard : std_logic;
	end record;
	constant init_digit : score_char := (score_rom_opcode => "0101010", score_top => 7, score_bottom => 23, score_left => 0, score_right => 0, fontBitEn => '0', inScoreboard => '0');--- ****** ---

	type type_scoreArray is array(natural range <>) of score_char;--- ****** ---


	----------------- SPECIAL ENEMY ROMs ----------------------

	type type_specialEnemy is array(natural range <>, natural range <>) of integer;

	constant specialEnemy15 : type_specialEnemy :=
	(
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,1,0,0,0,0,0,0,0,1,0,0,0),
		(0,0,0,0,1,0,0,0,0,0,1,0,0,0,0),
		(0,0,0,0,1,1,0,0,0,1,1,0,0,0,0),
		(0,0,0,1,1,1,1,1,1,1,1,1,0,0,0),
		(0,1,1,1,2,1,1,1,1,1,2,1,1,1,0),
		(0,1,1,1,1,1,1,1,1,1,1,1,1,1,0),
		(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
		(1,0,0,1,1,1,1,1,1,1,1,1,0,0,1),
		(1,0,0,1,0,0,0,0,0,0,0,1,0,0,1),
		(1,0,0,1,0,0,0,0,0,0,0,1,0,0,1),
		(0,0,0,0,1,1,1,0,1,1,1,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0)
	);

	constant specialEnemy25 : type_specialEnemy :=
	(
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
		(0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0),
		(0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0),
		(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
		(0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0),
		(0,0,1,1,1,1,1,2,2,1,1,1,1,1,1,1,2,2,1,1,1,1,1,0,0),
		(0,0,1,1,1,1,1,2,2,1,1,1,1,1,1,1,2,2,1,1,1,1,1,0,0),
		(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
		(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
		(1,1,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1),
		(1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,1,1),
		(1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1),
		(1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1),
		(1,1,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1),
		(0,0,0,0,0,0,0,1,1,1,1,0,0,1,1,1,1,1,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,1,1,1,1,0,0,1,1,1,1,1,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0)
	);

	constant specialEnemy30 : type_specialEnemy :=
	(
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0),
		(0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0),
		(0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
		(0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0),
		(0,0,0,1,1,1,1,1,2,2,2,1,1,1,1,1,1,1,1,2,2,2,1,1,1,1,1,0,0,0),
		(0,0,0,1,1,1,1,1,2,2,2,1,1,1,1,1,1,1,1,2,2,2,1,1,1,1,1,0,0,0),
		(0,0,0,1,1,1,1,1,2,2,2,1,1,1,1,1,1,1,1,2,2,2,1,1,1,1,1,0,0,0),
		(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
		(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
		(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
		(1,1,1,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1,1),
		(1,1,1,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1,1),
		(1,1,1,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1,1),
		(1,1,1,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,1,1,1),
		(1,1,1,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,1,1,1),
		(0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0)
	);

	------------ Alien ROMs -added by Nathan--

	type small_alien_rom_type is array (0 to 14) of std_logic_vector(0 to 14);
	constant small_alien_rom_const : small_alien_rom_type :=
	(
		"001100000001100",
		"000110000011100",
		"000111101111000",
		"000111111111000",
		"001111111111100",
		"011110111011110",
		"011111111111110",
		"010111111111010",
		"011111000111110",
		"010111111111010",
		"000011111110000",
		"000000000000000",
		"000000000000000",
		"000000000000000",
		"000000000000000"
	);

	type medium_alien_rom_type is array (0 to 24) of std_logic_vector(0 to 24);
	constant medium_alien_rom_const : medium_alien_rom_type :=
	(
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000011100000000011100000",
		"0000001100000000011000000",
		"0000000111000001110000000",
		"0000000111000001110000000",
		"0000011111111111111100000",
		"0000011111111111111100000",
		"0001111101111111011111000",
		"0001111101111111011111000",
		"0111111111111111111111110",
		"0111111111111111111111110",
		"0111011111111111111101110",
		"0111011111111111111101110",
		"0111011100000000011101110",
		"0010001100000000011000100",
		"0000000111110111110000000",
		"0000000011100011100000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000"
	);

	type large_alien_rom_type is array (0 to 29) of std_logic_vector(0 to 29);
	constant large_alien_rom_const : large_alien_rom_type :=
	(
		"000000000000000000000000000000",
		"000000000000000000000000000000",
		"000000011000000000000110000000",
		"000000011000000000000110000000",
		"000000011110000000011110000000",
		"000000000110000000011000000000",
		"000000000110000000011000000000",
		"000000011111111111111110000000",
		"000000011111111111111110000000",
		"000011111001111111100111110000",
		"000011111001111111100111110000",
		"000011111001111111100111110000",
		"001111111111111111111111111100",
		"001111111111111111111111111100",
		"001100011111111111111110001100",
		"001100011111111111111110001100",
		"001100011111111111111110001100",
		"001100011000000000000110001100",
		"001100011000000000000110001100",
		"000000000111110011111000000000",
		"000000000111110011111000000000",
		"000000000000000000000000000000",
		"000000000000000000000000000000",
		"000000000000000000000000000000",
		"000000000000000000000000000000",
		"000000000000000000000000000000",
		"000000000000000000000000000000",
		"000000000000000000000000000000",
		"000000000000000000000000000000",
		"000000000000000000000000000000"
	);


	signal alien_rom_addr , alien_rom_col : integer;
	signal alien_rom_data_15: std_logic_vector (0 to 14);
	signal alien_rom_data_25: std_logic_vector (0 to 24);
	signal alien_rom_data_30: std_logic_vector (0 to 29);
	signal alien_rom_bit : std_logic ;


	---------------------------- Object Roms --------------------------------------
	type object_rom_type is array (0 to 24) of std_logic_vector(0 to 24);
	constant met_object_rom_const : object_rom_type :=
	(
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000001001000000000000000",
		"0001111111111010000000000",
		"0011111111111110100000000",
		"0111111111111111111000000",
		"0111111111000111111111100",
		"1111111111010000111111110",
		"1111111111100011111111100",
		"0111111110011111111101000",
		"0011111111111111110000000",
		"0001111111111111100000000",
		"0000001111010000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000"
	);

	--type object_rom_type is array (0 to 24) of std_logic_vector(0 to 24);
	constant ufo_object_rom_const : object_rom_type :=
	(
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000001111100000000000",
		"0000000011111110000000000",
		"0000000011111110000000000",
		"0000000111111111100000000",
		"0001111111111111111100000",
		"0111111111111111100000110",
		"0000111111111111000000000",
		"0000000011111010000000000",
		"0000000001000010000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000"
	);

	--type object_rom_type is array (0 to 24) of std_logic_vector(0 to 24);
	constant sat_object_rom_const : object_rom_type :=
	(
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0111111111000001111111111",
		"1111111111101011111111111",
		"1111111111101011111111111",
		"0111111111111111111111111",
		"0000000000101110000000000",
		"0000000000101110000000000",
		"0000000000101110000000000",
		"0000000000101110000000000",
		"0000000000101110000000000",
		"0000000000001110000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000",
		"0000000000000000000000000"
	);



	-------------------------------------------------------------------------------


	-------------------------- SKY ------------------------------------------------

	type sky_data is
		record
			pixelOn : boolean;
			rgb : std_logic_vector(11 downto 0);
		end record;
	constant init_sky : sky_data := (pixelOn => false, rgb => "111111111111");

	-------------------------------------------------------------------------------

	---------------------------------------------------------------------------------------------------------------------------------------------------
	--RECORD TYPES:
	--Ship:
	constant init_ship_pos : point_2D := (x => shipsInitialx, y => shipsInitialy);
	constant init_ship_vel, init_enemy_vel: point_2D := (x => 0, y => 0);
	--Lasers:
	constant laser_velo : point_2D := (x => 25, y => 0);
	--Enemies:
	--Initalize to be off screen just in case
	constant smallPos : point_2D := (x => smallStartX, y => smallStartY);
	constant medPos : point_2D := (x => MedStartX, y => medStartY);
	constant bigPos : point_2D := (x => MedStartX, y => bigStartY);
	constant offScreen : point_2D := (x => 660, y => 500);
	constant small_Velo : point_2D :=(x => -5, y => 0);
	constant med_velo : point_2D := (x => -4, y => 0);
	constant big_velo : point_2D := (x => -3, y => 0);
	constant obj_velo : point_2D := (x=> objVeloX, y => objVeloY);
	constant obj_pos1 : point_2D := (x => objPosX, y => objPosy1);
	constant obj_pos2 : point_2D := (x => objPosX, y => objPosy2);
	constant obj_pos3 : point_2D := (x => objPosX, y => objPosy3);
	constant obj_pos4 : point_2D := (x => objPosX, y => objPosy4);
	constant obj_pos5 : point_2D := (x => objPosX, y => objPosy5);
	constant ZeroVelo : point_2D := (x => 0, y => 0);
	----------------------------------------------------------------------------------------------------------------------------------------------------
	type type_gameObj is
	record
		position : point_2D;
		ObjWidth : integer range 0 to 200;
		objHeight : integer range 0 to 200;
		velocity : point_2D;
		points : integer range 0 to 1000;
		element_on : boolean;
		lives : integer range 0 to 3;
		--lives
	end record;
	constant init_ship : type_gameObj    := (position => init_ship_pos, velocity => init_Ship_vel, objWidth => shipWidthConst, objHeight => shipHeightConst, points => 0, element_on => true, lives => 3);
	constant init_laser: type_gameObj    := (position => init_ship_pos, velocity => laser_velo, objWidth => laserWidth, objHeight => laserHeight, points => 0, element_on => false,lives => 0);

	constant init_small : type_gameObj   := (position => smallPos,   velocity => small_Velo,  objWidth => smallWidth, objHeight => smallHeight, points => 30, element_on => false,lives => 0);
	constant init_ShootingSmall : type_gameObj := (position => smallPos, velocity => small_Velo, objWidth => smallWidth, objHeight => smallHeight, points => 40, element_on => false, lives => 1);
	constant init_Med : type_gameObj     := (position => medPos ,    velocity => Med_Velo,    objWidth => medWidth,   objHeight => medHeight,   points => 18, element_on => false,lives => 0);
	constant init_ShootingMed : type_gameObj := (position => MedPos, velocity => Med_Velo, objWidth => MedWidth, objHeight => MedHeight, points => 30, element_on => false, lives => 1);
   constant init_Big : type_gameObj     := (position => bigPos ,    velocity => Big_Velo,    objWidth => bigWidth,   objHeight => bigHeight,   points => 10, element_on => false,lives => 0);
   constant init_ShootingBig : type_gameObj := (position => BigPos, velocity => Big_Velo, objWidth => BigWidth, objHeight => BigHeight, points => 30, element_on => false, lives => 1);
   constant zero_entries : type_gameObj := (position => offScreen,  velocity => ZeroVelo,     objWidth => 0,          objHeight => 0,           points => 0, element_on => false,lives => 0);

   constant init_obj1 : type_gameObj := (position => obj_pos1, velocity => obj_velo, objWidth => objectWidth, objHeight => objectHeight, points => 0, element_on => false, lives => 0);
    constant init_obj2 : type_gameObj := (position => obj_pos2, velocity => obj_velo, objWidth => objectWidth, objHeight => objectHeight, points => 0, element_on => false, lives => 0);
	constant init_obj3 : type_gameObj := (position => obj_pos3, velocity => obj_velo, objWidth => objectWidth, objHeight => objectHeight, points => 0, element_on => false, lives => 0);
  	constant init_obj4 : type_gameObj := (position => obj_pos4, velocity => obj_velo, objWidth => objectWidth, objHeight => objectHeight, points => 0, element_on => false, lives => 0);
	constant init_obj5 : type_gameObj := (position => obj_pos5, velocity => obj_velo, objWidth => objectWidth, objHeight => objectHeight, points => 0, element_on => false, lives => 0);
	--------------------------------------------------------------------------------------------------------------------------------------------------------------
	type type_gameObjArray is array(natural range <>) of type_gameObj;
	type type_gameObjMatrix is array(integer range 0 to 8, integer range 0 to 5) of type_gameObj;

   ------------------------------------------------------------------------------------------------------------------------------------------------------
	type type_bounds is
	record
		   L : integer range -8192 to 8191;
	      R : integer range -8192 to 8191;
	    top : integer range -8192 to 8191;
	 bottom : integer range -8192 to 8191;
	end record;
	--------------------------------------------------------------------------------------------------------
	type type_drawElement is
	record
		pixelOn : boolean;
		rgb : std_logic_vector(11 downto 0);
	end record;
	constant init_type_drawElement : type_drawElement := (pixelOn => false, rgb => (others => '0'));
	type drawElementArray is array(natural range <>) of type_drawElement;
	type drawElementMatrix is array(integer range 0 to 8, integer range 0 to 5) of type_drawElement;
	-------------------------------------------------------------------------------------------------------------------
	type controls is
	record
		up : std_logic;
		down: std_logic;
		L : std_logic;
		R : std_logic;
		moveMagx, moveMagy: std_logic_vector(2 downto 0);
		shoot : std_logic;
	end record;
	constant init_controls : controls := ('0','0','0','0',(others => '0'), (others => '0'), '0');
	------------------------------------------------------------------------
	-- Functions:
	function createBounds(object : type_gameobj) return type_Bounds;
	function checkCollisionX(obj1, obj2 : type_gameObj) return boolean;
	function checkCollisionY(obj1, obj2 : type_gameObj) return boolean;

end package graphicsPackage;
-----***********************************************************************************************************************************************

package body graphicsPackage is


	function createBounds(object : type_gameObj) return type_bounds is
		variable bounds : type_bounds;
	begin
		bounds.L := object.position.x;
		bounds.R := object.position.x + Object.objWidth-1;
		bounds.top := object.position.y;
		bounds.bottom := object.position.y + object.objHeight-1;
	return bounds;
   end function createbounds;

	function checkCollisionX(obj1, obj2 : type_gameObj) return boolean is
		variable obj1_bounds : type_bounds := createBounds(obj1);
		variable obj2_bounds : type_bounds := createBounds(obj2);
	begin
		return (obj1_bounds.R >= obj2_bounds.L AND obj1_bounds.R <= obj2_bounds.R)
			or (obj1_bounds.L >= obj2_bounds.L and obj1_bounds.L <= obj2_bounds.R);
  end checkCollisionX;

	function checkCollisionY(obj1, obj2 : type_gameObj) return boolean is
		variable obj1_bounds : type_bounds := createBounds(obj1);
		variable obj2_bounds : type_bounds := createBounds(obj2);
	begin
		return (obj1_bounds.top >= obj2_bounds.top AND obj1_bounds.top <= obj2_bounds.bottom)
			or (obj1_bounds.bottom >= obj2_bounds.top and obj1_bounds.bottom <= obj2_bounds.bottom);
  end checkCollisionY;
 ---------------------------------------------------------------------------------------------

end package body;
